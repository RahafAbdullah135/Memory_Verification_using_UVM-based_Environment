package pack ;
    `include "transaction.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "subscriber.sv"
    `include "scoreboard.sv"
    `include "env.sv"
endpackage